typedef enum bit [3:0] {PHASE_1, PHASE_2, PHASE_3} phases_t;

typedef enum bit [2:0] {D7, D6, D5, D4, D3, D2, D1, RW_, X} within_phase_t;