module OV7670_SIM (
    input clk,
    input reset,

    output logic hsync,
    output logic vsync,
    output logic [7:0] data,
    output logic pixclk
);

endmodule